module token

pub struct Pos {
pub:
	len     int
	pos     int
	col     int
}

