module ast

[heap]
pub struct Scope {
	start_pos int
	end_pos   int
}
