module main

import repl

fn main() {
	println('Monkey REPL')
	repl.start()
}
